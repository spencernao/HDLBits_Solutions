module top_module ( input a, input b, output out );
    mod_a instance1(.in2(b),.in1(a),.out(out));
endmodule
